module run();
  wire clk;
  clock c(clk);
  regbank_tb tb(clk);
endmodule